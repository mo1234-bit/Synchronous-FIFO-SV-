package shared_pkg;
	bit test_finished;
	int correct_count,errors_count;
endpackage : shared_pkg